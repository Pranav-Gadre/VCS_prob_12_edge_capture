module edge_capture (
	input   wire        clk,
	input   wire        reset,

	input   wire [31:0] data_i,

	output  wire [31:0] edge_o

);

	// Write your logic here...
	
	
endmodule